-- Hazards Unit 


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity forward_unit is
    port( instruction_in   : in std_logic_vector(15 downto 0);
          instruction_out : out std_logic_vector(15 downto 0)  
    );
  
end forward_unit;

architecture Behavioral of forward_unit is
  
  
  
  
  
  
end Behavioral;